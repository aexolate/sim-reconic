`timescale 1ns / 1ps

module s_axi_adapter_wrapper(
    input clk,
    input [7:0] s_axi_awid,
    input [63:0] s_axi_awaddr,
    input [7:0] s_axi_awlen,
    input [7:0] s_axi_awsize,
    input [2:0] s_axi_awburst,
    input s_axi_awvalid,
    output reg s_axi_awready,
    input [127:0] s_axi_wdata,
    input [15:0] s_axi_wstrb,
    input s_axi_wlast,
    input s_axi_wvalid,
    output reg s_axi_wready,
    output reg [7:0] s_axi_bid,
    output reg [1:0] s_axi_bresp,
    output reg s_axi_bvalid,
    input s_axi_bready,
    input [7:0] s_axi_arid,
    input [63:0] s_axi_araddr,
    input [7:0] s_axi_arlen,
    input [2:0] s_axi_arsize,
    input [2:0] s_axi_arburst,
    input s_axi_arvalid,
    output reg s_axi_arready,
    output reg [7:0] s_axi_rid,
    output reg [127:0] s_axi_rdata,
    output reg [1:0] s_axi_rresp,
    output reg s_axi_rlast,
    output reg s_axi_rvalid,
    input s_axi_rready
);

    s_axi_adapter s_axi_adapter_inst(
        .clk(clk),
        .s_axi_awid(s_axi_awid),
        .s_axi_awaddr(s_axi_awaddr),
        .s_axi_awlen(s_axi_awlen),
        .s_axi_awsize(s_axi_awsize),
        .s_axi_awburst(s_axi_awburst),
        .s_axi_awvalid(s_axi_awvalid),
        .s_axi_awready(s_axi_awready),
        .s_axi_wdata(s_axi_wdata),
        .s_axi_wstrb(s_axi_wstrb),
        .s_axi_wlast(s_axi_wlast),
        .s_axi_wvalid(s_axi_wvalid),
        .s_axi_wready(s_axi_wready),
        .s_axi_bid(s_axi_bid),
        .s_axi_bresp(s_axi_bresp),
        .s_axi_bvalid(s_axi_bvalid),
        .s_axi_bready(s_axi_bready),
        .s_axi_arid(s_axi_arid),
        .s_axi_araddr(s_axi_araddr),
        .s_axi_arlen(s_axi_arlen),
        .s_axi_arsize(s_axi_arsize),
        .s_axi_arburst(s_axi_arburst),
        .s_axi_arvalid(s_axi_arvalid),
        .s_axi_arready(s_axi_arready),
        .s_axi_rid(s_axi_rid),
        .s_axi_rdata(s_axi_rdata),
        .s_axi_rresp(s_axi_rresp),
        .s_axi_rlast(s_axi_rlast),
        .s_axi_rvalid(s_axi_rvalid),
        .s_axi_rready(s_axi_rready)
    );
    
endmodule